module timer();


 